`ifndef __FUNCTIONS__
`define __FUNCTIONS__

module functions;

endmodule


`endif