module ParallelImageProcessor #(
) (
);


endmodule;